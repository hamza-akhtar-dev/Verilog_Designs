//------------------------------------------------------------------
// 			 Datapath for Unsigned Binary Multiplier
//------------------------------------------------------------------
module Datapath(
input[2:0] inA, inB,
input clk, loadRegs, addRegs, shiftReg, decrement,
output Zbit, Mbit,
output[5:0] product
);

reg [2:0] A, B, Q;
reg [1:0] P;
reg C;

always @ (posedge clk) 
begin

//------------------------------------------------------------------
//                      LOADING REGISTERS    
//------------------------------------------------------------------

if (loadRegs) 
begin
	P <= 3;
	A <= 0;
	C <= 0;
	B <= inA;
	Q <= inB;
end

//------------------------------------------------------------------
//                            ADDER
//------------------------------------------------------------------
if (addRegs) 
	{C, A} <= A + B;
	
//------------------------------------------------------------------
//                        SHIFT REGISTER
//------------------------------------------------------------------
if (shiftReg) 
	{C, A, Q} <= {C, A, Q} >> 1;
	
//------------------------------------------------------------------
//                        DOWN COUNTER
//------------------------------------------------------------------
if (decrement) 
	P <= P - 1;
end

assign Zbit = (P == 0);
assign Mbit = Q[0];
assign product = {A, Q};

endmodule